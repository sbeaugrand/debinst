.title KiCad schematic
R1 Net-_C17-Pad1_ Net-_J1-Pad1_ <R1>
C17 Net-_C17-Pad1_ GND <C17>
C18 sortie GND <C18>
R2 sortie GND <R2>
L4 Net-_C17-Pad1_ sortie <L4>
VJ1 Net-_J1-Pad1_ GND dc 0 ac <VJ1>
.control
ac dec 100 2Meg 8Meg
run
wrdata build/<dst> db(abs(V(sortie)))
.endc
.end
